* The classic RC filter!
V1 inp 0 DC 0 SIN(0 1 1k)
R1 inp out 1
C2 out 0 0.1m
.tran 1u 2m
.END